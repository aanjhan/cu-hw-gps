// megafunction wizard: %LPM_MULT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mult 

// ============================================================
// File Name: multiplier.v
// Megafunction Name(s):
// 			lpm_mult
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 8.0 Build 215 05/29/2008 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2008 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module dll_multiplier (
    input                          clock,
    input [INPUT_A_WIDTH-1:0]      dataa,
    input [INPUT_B_WIDTH-1:0]      datab,
    output wire [OUTPUT_WIDTH-1:0] result);

   parameter INPUT_A_WIDTH = 9;
   parameter INPUT_B_WIDTH = 9;
   parameter OUTPUT_WIDTH = 18;

   wire [OUTPUT_WIDTH-1:0] sub_wire0;
   assign result = sub_wire0;

   lpm_mult lpm_mult_component (.dataa (dataa),
				.datab (datab),
				.clock (clock),
				.result (sub_wire0),
				.aclr (1'b0),
				.clken (1'b1),
				.sum (1'b0));
   defparam lpm_mult_component.lpm_hint = "MAXIMIZE_SPEED=9",
	    lpm_mult_component.lpm_pipeline = 2,
	    lpm_mult_component.lpm_representation = "UNSIGNED",
	    lpm_mult_component.lpm_type = "LPM_MULT",
	    lpm_mult_component.lpm_widtha = INPUT_A_WIDTH,
	    lpm_mult_component.lpm_widthb = INPUT_B_WIDTH,
	    lpm_mult_component.lpm_widthp = OUTPUT_WIDTH;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
// Retrieval info: PRIVATE: ConstantB NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "2"
// Retrieval info: PRIVATE: Latency NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
// Retrieval info: PRIVATE: SignedMult NUMERIC "0"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "1"
// Retrieval info: PRIVATE: WidthA NUMERIC "8"
// Retrieval info: PRIVATE: WidthB NUMERIC "8"
// Retrieval info: PRIVATE: WidthP NUMERIC "16"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: optimize NUMERIC "1"
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=9"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "2"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
// Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "8"
// Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "8"
// Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "16"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: dataa 0 0 8 0 INPUT NODEFVAL dataa[7..0]
// Retrieval info: USED_PORT: datab 0 0 8 0 INPUT NODEFVAL datab[7..0]
// Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT NODEFVAL result[15..0]
// Retrieval info: CONNECT: @dataa 0 0 8 0 dataa 0 0 8 0
// Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
// Retrieval info: CONNECT: @datab 0 0 8 0 datab 0 0 8 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier_bb.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier_waveforms.html FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier_wave*.jpg FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL multiplier_syn.v TRUE
// Retrieval info: LIB_FILE: lpm
