// This file is part of the Cornell University Hardware GPS Receiver Project.
// Copyright (C) 2009 - Adam Shapiro (ams348@cornell.edu)
//                      Tom Chatt (tjc42@cornell.edu)
//
// This program is free software; you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation; either version 2 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA

//This file was automatically generated by
//Matlab on 31-May-2009 12:11:08.
`include "sin.vh"

module sin(
    input [`SIN_INPUT_RANGE]       in,
    output reg [`SIN_OUTPUT_RANGE] out);

   always @(in) begin
     casez(in)
       `SIN_INPUT_WIDTH'd0: out <= `SIN_OUTPUT_WIDTH'd0;
       `SIN_INPUT_WIDTH'd1: out <= `SIN_OUTPUT_WIDTH'd1;
       `SIN_INPUT_WIDTH'd2: out <= `SIN_OUTPUT_WIDTH'd2;
       `SIN_INPUT_WIDTH'd3: out <= `SIN_OUTPUT_WIDTH'd3;
       `SIN_INPUT_WIDTH'd4: out <= `SIN_OUTPUT_WIDTH'd3;
       `SIN_INPUT_WIDTH'd5: out <= `SIN_OUTPUT_WIDTH'd3;
       `SIN_INPUT_WIDTH'd6: out <= `SIN_OUTPUT_WIDTH'd2;
       `SIN_INPUT_WIDTH'd7: out <= `SIN_OUTPUT_WIDTH'd1;
       `SIN_INPUT_WIDTH'd8: out <= `SIN_OUTPUT_WIDTH'd5;
       `SIN_INPUT_WIDTH'd9: out <= `SIN_OUTPUT_WIDTH'd6;
       `SIN_INPUT_WIDTH'd10: out <= `SIN_OUTPUT_WIDTH'd7;
       `SIN_INPUT_WIDTH'd11: out <= `SIN_OUTPUT_WIDTH'd7;
       `SIN_INPUT_WIDTH'd12: out <= `SIN_OUTPUT_WIDTH'd7;
       `SIN_INPUT_WIDTH'd13: out <= `SIN_OUTPUT_WIDTH'd6;
       `SIN_INPUT_WIDTH'd14: out <= `SIN_OUTPUT_WIDTH'd5;
       `SIN_INPUT_WIDTH'd15: out <= `SIN_OUTPUT_WIDTH'd0;
       default: out <= `SIN_OUTPUT_WIDTH'hx;
     endcase
   end
endmodule
